// Belinda Brown Ramírez
// Brandon Esquivel Molina
// December, 2020
// timna.brown@ucr.ac.cr
// brandon.esquivel@ucr.ac.cr
//github: @brown9804, @brandonEsquivel

`timescale 1 ns / 1 ps

module system (
	input            clk,
	input            resetn,
	input 			 PS2Clk,
	input 			 PS2Data,
	output           trap,
	output reg [7:0] out_byte,
	output reg       out_byte_en,
	output reg [7:0] Anode_on,
    output reg [7:0] Led_output
);
	// set this to 0 for better timing but less performance/MHz
	parameter FAST_MEMORY = 1;

	// 4096 32bit words = 16kB memory
	parameter MEM_SIZE = 4096;

	wire mem_valid;
	wire mem_instr;
	reg mem_ready;
	wire [31:0] mem_addr;
	wire [31:0] mem_wdata;
	wire [3:0] mem_wstrb;
	reg [31:0] mem_rdata;

	wire mem_la_read;
	wire mem_la_write;
	wire [31:0] mem_la_addr;
	wire [31:0] mem_la_wdata;
	wire [3:0] mem_la_wstrb;

	picorv32 picorv32_core (
		.clk         (clk         ),
		.resetn      (resetn      ),
		.trap        (trap        ),
		.mem_valid   (mem_valid   ),
		.mem_instr   (mem_instr   ),
		.mem_ready   (mem_ready   ),
		.mem_addr    (mem_addr    ),
		.mem_wdata   (mem_wdata   ),
		.mem_wstrb   (mem_wstrb   ),
		.mem_rdata   (mem_rdata   ),
		.mem_la_read (mem_la_read ),
		.mem_la_write(mem_la_write),
		.mem_la_addr (mem_la_addr ),
		.mem_la_wdata(mem_la_wdata),
		.mem_la_wstrb(mem_la_wstrb)
	);
	
// ------------------------------------------
// ////// -> BEGIN LAB8
// //////// begin part1
// text_display text_display_inst(
// // INPUTS 
// .clk (clk),
// .resetn (resetn),
// .select (out_byte[3:0]), // 4 bits // selector 
// .enable (out_byte_en), // 1 bit 
// // OUTPUTS
// .catode ( wled  ), // 7 segments 
// .anode (  wanode )
// );

///////// begin part2

prs_game  prs_game_inst(
// INPUTS 
.clk (clk),
.resetn (resetn),
.PS2Clk (PS2Clk),
.PS2Data (PS2Data),
// OUTPUTS
.catode ( wled  ), // 7 segments 
.anode (  wanode )
);
////// -> END LAB8
// ------------------------------------------
reg [31:0] memory [0:MEM_SIZE-1];

`ifdef SYNTHESIS
    initial $readmemh("../firmware/firmware.hex", memory);
`else
	initial $readmemh("firmware.hex", memory);
`endif

reg [31:0] m_read_data;
reg m_read_en;

generate if (FAST_MEMORY) begin
	always @(posedge clk) begin
		mem_ready <= 1;
		out_byte_en <= 0;
		mem_rdata <= memory[mem_la_addr >> 2];
		if (mem_la_write && (mem_la_addr >> 2) < MEM_SIZE) begin
			if (mem_la_wstrb[0]) memory[mem_la_addr >> 2][ 7: 0] <= mem_la_wdata[ 7: 0];
			if (mem_la_wstrb[1]) memory[mem_la_addr >> 2][15: 8] <= mem_la_wdata[15: 8];
			if (mem_la_wstrb[2]) memory[mem_la_addr >> 2][23:16] <= mem_la_wdata[23:16];
			if (mem_la_wstrb[3]) memory[mem_la_addr >> 2][31:24] <= mem_la_wdata[31:24];
		end
		else
		if (mem_la_write && mem_la_addr == 32'h1000_0000) begin
			out_byte_en <= 1;
			out_byte <= mem_la_wdata;
		end
	end
	end 
	else begin
		always @(posedge clk) begin
			m_read_en <= 0;
			mem_ready <= mem_valid && !mem_ready && m_read_en;

			m_read_data <= memory[mem_addr >> 2];
			mem_rdata <= m_read_data;

			out_byte_en <= 0;

			(* parallel_case *)
			case (1)
				mem_valid && !mem_ready && !mem_wstrb && (mem_addr >> 2) < MEM_SIZE: begin
					m_read_en <= 1;
				end
				mem_valid && !mem_ready && |mem_wstrb && (mem_addr >> 2) < MEM_SIZE: begin
					if (mem_wstrb[0]) memory[mem_addr >> 2][ 7: 0] <= mem_wdata[ 7: 0];
					if (mem_wstrb[1]) memory[mem_addr >> 2][15: 8] <= mem_wdata[15: 8];
					if (mem_wstrb[2]) memory[mem_addr >> 2][23:16] <= mem_wdata[23:16];
					if (mem_wstrb[3]) memory[mem_addr >> 2][31:24] <= mem_wdata[31:24];
					mem_ready <= 1;
				end
				mem_valid && !mem_ready && |mem_wstrb && mem_addr == 32'h1000_0000: begin
					out_byte_en <= 1;
					out_byte <= mem_wdata;
					mem_ready <= 1;
				end
			endcase
		end
	end 
endgenerate


//// Exe 1 wires ///
wire [7:0] wanode;
wire [7:0] wled;

/////// Logic /////////////////////
	always @(posedge clk) begin
	   if (~resetn) begin
	       Anode_on         <= 8'b11111111;
	       Led_output       <= 8'b11111111;
	   end 
	   else begin
           Anode_on        <= wanode;
	       Led_output      <= wled;
	   end
	end

/////////////////////////////////

endmodule
